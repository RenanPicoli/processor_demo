mem_code_for_7seg_inst : mem_code_for_7seg PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
